`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.06.2025 17:17:42
// Design Name: 
// Module Name: tb_mux2to1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps

module tb_mux2to1;

    reg a, b, sel;
    wire y;

    mux2to1 uut (
        .a(a),
        .b(b),
        .sel(sel),
        .y(y)
    );

    initial begin
        a = 0; b = 1; sel = 0;
        #10 sel = 1;
        #10 a = 1; b = 0; sel = 0;
        #10 sel = 1;
        #10 $finish;
    end

    initial begin
        $monitor("Time=%0t | a=%b b=%b sel=%b => y=%b", $time, a, b, sel, y);
    end

endmodule
